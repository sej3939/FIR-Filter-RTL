
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   sj3939@hansolo.poly.edu
//  Generated date: Thu Dec 12 20:33:31 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output, Shift_Accum_Loop_C_6_tr0
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input Shift_Accum_Loop_C_6_tr0;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    Shift_Accum_Loop_C_0 = 4'd1,
    Shift_Accum_Loop_C_1 = 4'd2,
    Shift_Accum_Loop_C_2 = 4'd3,
    Shift_Accum_Loop_C_3 = 4'd4,
    Shift_Accum_Loop_C_4 = 4'd5,
    Shift_Accum_Loop_C_5 = 4'd6,
    Shift_Accum_Loop_C_6 = 4'd7,
    main_C_1 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      Shift_Accum_Loop_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = Shift_Accum_Loop_C_1;
      end
      Shift_Accum_Loop_C_1 : begin
        fsm_output = 9'b000000100;
        state_var_NS = Shift_Accum_Loop_C_2;
      end
      Shift_Accum_Loop_C_2 : begin
        fsm_output = 9'b000001000;
        state_var_NS = Shift_Accum_Loop_C_3;
      end
      Shift_Accum_Loop_C_3 : begin
        fsm_output = 9'b000010000;
        state_var_NS = Shift_Accum_Loop_C_4;
      end
      Shift_Accum_Loop_C_4 : begin
        fsm_output = 9'b000100000;
        state_var_NS = Shift_Accum_Loop_C_5;
      end
      Shift_Accum_Loop_C_5 : begin
        fsm_output = 9'b001000000;
        state_var_NS = Shift_Accum_Loop_C_6;
      end
      Shift_Accum_Loop_C_6 : begin
        fsm_output = 9'b010000000;
        if ( Shift_Accum_Loop_C_6_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = Shift_Accum_Loop_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b100000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = Shift_Accum_Loop_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, y_rsc_dat, y_triosy_lz, x_rsc_dat, x_triosy_lz
);
  input clk;
  input rst;
  output [7:0] y_rsc_dat;
  output y_triosy_lz;
  input [7:0] x_rsc_dat;
  output x_triosy_lz;


  // Interconnect Declarations
  wire [7:0] x_rsci_idat;
  reg [6:0] y_rsci_idat_7_1;
  reg y_rsci_idat_0;
  wire [8:0] fsm_output;
  wire [3:0] Shift_Accum_Loop_acc_1_tmp;
  wire [4:0] nl_Shift_Accum_Loop_acc_1_tmp;
  wire and_dcpl_1;
  wire or_dcpl_10;
  wire or_tmp_3;
  wire or_tmp_19;
  wire and_21_cse;
  reg [2:0] i_3_0_sva_2_0;
  reg i_3_0_sva_1_3;
  reg reg_x_triosy_obj_ld_cse;
  wire or_tmp_23;
  wire [7:0] z_out;
  wire [8:0] nl_z_out;
  reg [7:0] shift_reg_0_lpi_2;
  reg [7:0] shift_reg_2_lpi_2;
  reg [7:0] shift_reg_3_lpi_2;
  reg [7:0] shift_reg_1_lpi_2;
  reg [7:0] shift_reg_4_lpi_2;
  reg [7:0] x_sva;
  reg [6:0] acc_sva_7_1;
  reg acc_sva_0;
  wire [7:0] Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1;
  wire [2:0] Shift_Accum_Loop_else_acc_1_tmp;
  wire [3:0] nl_Shift_Accum_Loop_else_acc_1_tmp;
  wire [7:0] Shift_Accum_Loop_else_mul_itm;
  wire [10:0] nl_Shift_Accum_Loop_else_mul_itm;

  wire[6:0] mux_nl;
  wire acc_not_nl;
  wire Shift_Accum_Loop_mux_4_nl;
  wire or_27_nl;
  wire[2:0] Shift_Accum_Loop_else_mux_5_nl;
  wire Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_2_nl;
  wire[5:0] Shift_Accum_Loop_if_mux_4_nl;
  wire Shift_Accum_Loop_if_mux_5_nl;
  wire Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_3_nl;
  wire[6:0] Shift_Accum_Loop_if_mux_6_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_y_rsci_idat;
  assign nl_y_rsci_idat = {y_rsci_idat_7_1 , y_rsci_idat_0};
  ccs_out_v1 #(.rscid(32'sd1),
  .width(32'sd8)) y_rsci (
      .idat(nl_y_rsci_idat[7:0]),
      .dat(y_rsc_dat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd8)) x_rsci (
      .dat(x_rsc_dat),
      .idat(x_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) y_triosy_obj (
      .ld(reg_x_triosy_obj_ld_cse),
      .lz(y_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) x_triosy_obj (
      .ld(reg_x_triosy_obj_ld_cse),
      .lz(x_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .Shift_Accum_Loop_C_6_tr0(i_3_0_sva_1_3)
    );
  assign nl_Shift_Accum_Loop_else_acc_1_tmp = i_3_0_sva_2_0 + 3'b111;
  assign Shift_Accum_Loop_else_acc_1_tmp = nl_Shift_Accum_Loop_else_acc_1_tmp[2:0];
  assign Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1
      = MUX_v_8_5_2(shift_reg_0_lpi_2, shift_reg_1_lpi_2, shift_reg_2_lpi_2, shift_reg_3_lpi_2,
      shift_reg_4_lpi_2, Shift_Accum_Loop_else_acc_1_tmp);
  assign nl_Shift_Accum_Loop_acc_1_tmp = conv_u2s_3_4(i_3_0_sva_2_0) + 4'b1111;
  assign Shift_Accum_Loop_acc_1_tmp = nl_Shift_Accum_Loop_acc_1_tmp[3:0];
  assign and_dcpl_1 = ~((fsm_output[8]) | (fsm_output[0]));
  assign or_dcpl_10 = (i_3_0_sva_2_0!=3'b000);
  assign or_tmp_3 = (fsm_output[8]) | (fsm_output[0]);
  assign and_21_cse = (i_3_0_sva_2_0==3'b000) & (fsm_output[1]);
  assign or_tmp_19 = ~(i_3_0_sva_1_3 & (fsm_output[7]));
  assign or_tmp_23 = or_dcpl_10 & (fsm_output[1]);
  assign Shift_Accum_Loop_else_mux_5_nl = MUX_v_3_6_2x0(3'b000, 3'b101, 3'b101, 3'b000,
      3'b010, i_3_0_sva_2_0);
  assign nl_Shift_Accum_Loop_else_mul_itm = Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1
      * Shift_Accum_Loop_else_mux_5_nl;
  assign Shift_Accum_Loop_else_mul_itm = nl_Shift_Accum_Loop_else_mul_itm[7:0];
  always @(posedge clk) begin
    if ( rst ) begin
      acc_sva_7_1 <= 7'b0000000;
    end
    else if ( (fsm_output[0]) | (fsm_output[8]) | (fsm_output[1]) ) begin
      acc_sva_7_1 <= MUX_v_7_2_2(7'b0000000, mux_nl, acc_not_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_sva <= 8'b00000000;
    end
    else if ( ~ and_dcpl_1 ) begin
      x_sva <= x_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      acc_sva_0 <= 1'b0;
      reg_x_triosy_obj_ld_cse <= 1'b0;
    end
    else begin
      acc_sva_0 <= Shift_Accum_Loop_mux_4_nl & (~ or_tmp_3);
      reg_x_triosy_obj_ld_cse <= i_3_0_sva_1_3 & (fsm_output[7]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_3_0_sva_2_0 <= 3'b000;
    end
    else if ( or_tmp_3 | (fsm_output[1]) ) begin
      i_3_0_sva_2_0 <= MUX_v_3_2_2(3'b101, (Shift_Accum_Loop_acc_1_tmp[2:0]), fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_0_lpi_2 <= 8'b00000000;
    end
    else if ( (~ or_dcpl_10) & (fsm_output[1]) ) begin
      shift_reg_0_lpi_2 <= x_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_1_lpi_2 <= 8'b00000000;
    end
    else if ( (i_3_0_sva_2_0[0]) & (~ (i_3_0_sva_2_0[2])) & (fsm_output[1]) & (~
        (i_3_0_sva_2_0[1])) & ((Shift_Accum_Loop_else_acc_1_tmp!=3'b001)) ) begin
      shift_reg_1_lpi_2 <= Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_2_lpi_2 <= 8'b00000000;
    end
    else if ( (~((i_3_0_sva_2_0[0]) | (i_3_0_sva_2_0[2]))) & (fsm_output[1]) & (i_3_0_sva_2_0[1])
        & ((Shift_Accum_Loop_else_acc_1_tmp!=3'b010)) ) begin
      shift_reg_2_lpi_2 <= Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_3_lpi_2 <= 8'b00000000;
    end
    else if ( (i_3_0_sva_2_0[0]) & (~ (i_3_0_sva_2_0[2])) & (fsm_output[1]) & (i_3_0_sva_2_0[1])
        & ((Shift_Accum_Loop_else_acc_1_tmp!=3'b011)) ) begin
      shift_reg_3_lpi_2 <= Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_4_lpi_2 <= 8'b00000000;
    end
    else if ( (i_3_0_sva_2_0==3'b100) & (fsm_output[1]) & ((Shift_Accum_Loop_else_acc_1_tmp!=3'b100))
        ) begin
      shift_reg_4_lpi_2 <= Shift_Accum_Loop_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_0 <= 1'b0;
    end
    else if ( ~ or_tmp_19 ) begin
      y_rsci_idat_0 <= acc_sva_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_7_1 <= 7'b0000000;
    end
    else if ( ~ or_tmp_19 ) begin
      y_rsci_idat_7_1 <= acc_sva_7_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_3_0_sva_1_3 <= 1'b0;
    end
    else if ( fsm_output[1] ) begin
      i_3_0_sva_1_3 <= Shift_Accum_Loop_acc_1_tmp[3];
    end
  end
  assign mux_nl = MUX_v_7_2_2((z_out[7:1]), (z_out[6:0]), and_21_cse);
  assign acc_not_nl = ~ or_tmp_3;
  assign or_27_nl = (and_dcpl_1 & (~ (fsm_output[1]))) | and_21_cse;
  assign Shift_Accum_Loop_mux_4_nl = MUX_s_1_2_2((z_out[0]), acc_sva_0, or_27_nl);
  assign Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_2_nl = (acc_sva_7_1[6]) & or_tmp_23;
  assign Shift_Accum_Loop_if_mux_4_nl = MUX_v_6_2_2((acc_sva_7_1[6:1]), (acc_sva_7_1[5:0]),
      or_tmp_23);
  assign Shift_Accum_Loop_if_mux_5_nl = MUX_s_1_2_2((acc_sva_7_1[0]), acc_sva_0,
      or_tmp_23);
  assign Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_3_nl = (Shift_Accum_Loop_else_mul_itm[7])
      & or_tmp_23;
  assign Shift_Accum_Loop_if_mux_6_nl = MUX_v_7_2_2((x_sva[6:0]), (Shift_Accum_Loop_else_mul_itm[6:0]),
      or_tmp_23);
  assign nl_z_out = ({Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_2_nl , Shift_Accum_Loop_if_mux_4_nl
      , Shift_Accum_Loop_if_mux_5_nl}) + ({Shift_Accum_Loop_if_Shift_Accum_Loop_if_and_3_nl
      , Shift_Accum_Loop_if_mux_6_nl});
  assign z_out = nl_z_out[7:0];

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_6_2x0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      default : begin
        result = input_5;
      end
    endcase
    MUX_v_3_6_2x0 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_5_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      default : begin
        result = input_4;
      end
    endcase
    MUX_v_8_5_2 = result;
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tt_um_fir
// ------------------------------------------------------------------


module tt_um_fir (
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(~rst_n),
      .y_rsc_dat(uo_out),
    .y_triosy_lz(),
      .x_rsc_dat(ui_in),
    .x_triosy_lz()
    );
  assign uio_out = 8'b00000000;
  assign uio_oe = 8'b00000000;
endmodule



